/////////data flow ////////
module mux81 (input [7:0]I,
              input [2:0]s,
              output y);
assign y =((~s[0]) & (~s[1]) & (~s[2]) & I[0]) | 
           ((~s[0]) & (~s[1]) & (s[2]) & I[1]) | 
           ((~s[0]) & (s[1]) & (~s[2]) & I[2]) | 
           ((~s[0]) & (s[1]) & (s[2]) & I[3]) | 
           ((s[0]) & (~s[1]) & (~s[2]) & I[4]) | 
           ((s[0]) & (~s[1]) & (s[2]) & I[5]) | 
           ((s[0]) & (s[1]) & (~s[2]) & I[6]) | 
           ((s[0]) & (s[1]) & (s[2]) & I[7]);
endmodule           
